//                      FFT32_original                   //
// NO PIPELINE, only insert register in input and output. //



module FFT32_original (
		input clk,
		input i_rst,
		?
);

? 
endmodule




